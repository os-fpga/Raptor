module logic0 (logic0);
output logic0;
wire logic0;
assign logic0 = 1'b0;
endmodule
