`timescale 1 ps/ 1 ps 
///////////////////////////////////////////////////////////////// 
// Company: 
// Engineer: 
// Create Date: 2022-07-01 16:34:14
// Design Name: 
// Module Name: use_ip
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision: 
// Additional Comments:
// 
///////////////////////////////////////////////////////////////// 


module use_ip( 

    ); 
endmodule 
