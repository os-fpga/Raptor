module const1
(
    const1
);

    output const1;

    wire const1;

    TIEHBWP7D5T16P96CPD tiehi_U1 (.Z(const1));


endmodule

