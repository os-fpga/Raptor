module const0
(
    const0
);

    output const0;

    wire const0;

    TIELBWP7D5T16P96CPD tielo_U1 (.ZN(const0));

endmodule

