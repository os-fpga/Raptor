module bottom (input logic [`P1:0] a, output logic [`P1:0] b);
assign b = a;
endmodule
