module inverter (a,z);
input a;
output z;
wire z;
//assign z = ~a;
INVD4BWP7D5T16P96CPD U0 (.I(a), .ZN(z));
endmodule
