`include "def.vh"
module top(input logic [`P2:0] a, output logic [`P2:0] b);
   bottom bot (a, b);
   
   
endmodule // top

