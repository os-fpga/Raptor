`timescale 1 ps/ 1 ps 
////////////////////////////////////////////////////////////////////////////////// 
// Company: 
// Engineer: 
// Create Date: 2021-12-03 18:02:58
// Design Name: 
// Module Name: test
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision: 
// Additional Comments:
// 
////////////////////////////////////////////////////////////////////////////////// 


module test( 

    ); 
endmodule 
