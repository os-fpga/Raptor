`ifndef BRAM_SV_H
`define BRAM_SV_H
   localparam MODE_36  = 3'b011;  //36 or 32-bit 
   localparam MODE_18  = 3'b010; // 18 or  16-bit 
   localparam MODE_9   = 3'b001;   // 9 or 8-bit  
   localparam MODE_4   = 3'b100;   // 4-bit
   localparam MODE_2   = 3'b110; //32-bit
   localparam MODE_1   = 3'b101; //32-bit
`endif
