module logic1
(
    logic1
);

    output logic1;

    wire logic1;

    TIEHBWP7D5T16P96CPD tiehi_U1 (.Z(logic1));


endmodule

