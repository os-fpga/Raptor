module logic1 (logic1);
output logic1;
wire logic1;
assign logic1 = 1'b1;
endmodule
