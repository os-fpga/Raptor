module logic0
(
    logic0
);

    output logic0;

    wire logic0;

    TIELBWP7D5T16P96CPD tielo_U1 (.ZN(logic0));

endmodule

